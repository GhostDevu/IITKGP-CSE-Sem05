`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Computer Organization Laboratory (CS39001)
// Semester 05 (Autumn 2021-22)
// Assignment 06 -- Problem 02 [Bit Serial Adder]
// 		File Summary : Designed and implemented a Bit Serial Adder
// Group No. 16
//      Hritaban Ghosh (19CS30053)
//      Nakul Aggarwal (19CS10044)
//////////////////////////////////////////////////////////////////////////////////
// [[ Bit Serial Adder ]] -- Module for Bit Serial Adder (takes in three 1- bit inputs
// 'clk', 'rst' and 'load' and two 8-bit inputs 'input_A' and 'input_B' and outputs one
// 8-bit output 'sum' and one 1-bit output 'carry_out'.
//////////////////////////////////////////////////////////////////////////////////
// The 8-Bit Serial Adder circuit, which can perform addition in just 8 clock cycles.
//////////////////////////////////////////////////////////////////////////////////
module Bit_Serial_Adder(clk, rst, load, carry_out, sum, input_A, input_B);
	input wire [7:0] input_A, input_B;		// input_A and input_B are the operands of the addition operation
	input wire clk, rst, load;		// clk is the clock signal, rst is the reset signal and load is the signal to indicate that inputs are to be loaded
	output wire [7:0] sum;			// sum outputs the addition sum of input_A and input_B
	output reg carry_out;			// carry_out outputs the last carry_out of the addition process
	
	// Interconnecting Wires
	// a - 1-bit input from A
	// b - 1-bit input from B
	// s - sum of a and b
	// cout - carry out bit generated when a and b are added
	// cin - carry in bit from the previous addition
	wire a, b, s, cout, cin; 
	
	// Two Input Parallel In Serial Out Right Shift Registers to hold input_A and input_B and keep spitting LSBs from the right
	PISO_Right_Shift_Register_8_bit R1( .clk(clk) , .rst(rst) , .load(load) , .inp(input_A) , .data(a)) ;
	PISO_Right_Shift_Register_8_bit R2( .clk(clk) , .rst(rst) , .load(load) , .inp(input_B) , .data(b)) ;
	
	// One Output Serial In Parallel Out Right Shift Registers which stores the sum of input_A and input_B and gives it as output
	SIPO_Right_Shift_Register_8_bit S( .clk(clk) , .rst(rst) , .load(load) , .inp(8'b00000000) , .fill_bit(s), .out(sum)) ;
	
	// One Full Adder Module to Perform Serial Addition
	Full_Adder FA( .a(a) , .b(b) , .carry_in(cin) , .sum(s) , .carry_out(cout));
	
	// One D-Flip Flop to store the carry out bit generated by the FA from the previous clock cycle to give it as input to the FA in the current clock cycle
	D_Flip_Flop DFF( .clk(clk), .rst(rst), .D(cout), .Q(cin));
	
	always @ (*)
		carry_out = cin; // The last carry generated as input for the full adder is the carry out bit of the whole addition
endmodule
